module RegBank
#(parameter WIDTH = 4, SIZE = 3)
(
 input            clk,
 input            we3,
 input [SIZE-1:0] A1,
 input [SIZE-1:0] A2,
 input [SIZE-1:0] A3,
 input [WIDTH-1:0] WD3,
 output [WIDTH-1:0] RD1,
 output [WIDTH-1:0] RD2
);

endmodule
