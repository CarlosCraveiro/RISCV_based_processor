module register
#( parameter WIDTH = 1 )
   (
    input  clk,
    input  in_data,
    input  enable,
    output ou_data
    );

endmodule
